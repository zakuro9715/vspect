module ui

fn test_divider() {
	assert divider('-', 10) == '----------'
}
